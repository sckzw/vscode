module SAMPLE(
    input CLK,
    input RSTX,
    input PSEL,
    input PENABLE,
    input [31:0] PADDR,
    input PWRITE,
    input [3:0] PSTRB,
    input [31:0] PWDATA,
    output PREADY,
    output [31:0] PRDATA,
);


    reg aaa;



endmodule

